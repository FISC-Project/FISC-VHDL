LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.numeric_std.all;
USE IEEE.std_logic_unsigned.all;
USE work.FISC_DEFINES.all;

ENTITY ALU IS
	PORT(
		clk    : in  std_logic;
		opA    : in  std_logic_vector(FISC_INTEGER_SZ-1 downto 0);
		opB    : in  std_logic_vector(FISC_INTEGER_SZ-1 downto 0);
		func   : in  std_logic_vector(3 downto 0);
		zero   : out std_logic;
		result : out std_logic_vector(FISC_INTEGER_SZ-1 downto 0)
	);
END;

ARCHITECTURE RTL OF ALU IS
	signal result_reg : std_logic_vector(FISC_INTEGER_SZ-1 downto 0) := (others => '0');
BEGIN
	result_reg <= 
		opA and opB WHEN func = "0000" ELSE -- AND
		opA or opB  WHEN func = "0001" ELSE -- ORR
		opA + opB   WHEN func = "0010" ELSE -- ADD
		opA - opB   WHEN func = "0110" ELSE -- SUB
		opB         WHEN func = "0111" ELSE -- pass operand B
		not (opA or opB) WHEN func =  "1100"; -- NOR

	result <= result_reg;
	zero   <= '1' WHEN result_reg = (result_reg'range => '0') ELSE '0';
END ARCHITECTURE RTL;